Non Inverting Amplifier:

* Created on 21 March 2018
* @author: Omama Elrefaei

* Accessing subcircuit:
Xopamp 1 2 3 opamp
* Signal source::
Vin 2 0 DC 1
*Vin 2 0 AC 1
* Circuit componants:
*.PARAM Rf = 1
R 3 0 1K
Rf 3 1 9K
* Analysis request:
.TF V(1) Vin
*.STEP PARAM Rf LIST 9k 19k
*.AC DEC 100 100 100G
* Subcircuit
.SUBCKT opamp 1 	2   	3
* Connection: | 	|  		|
*   		o/p 	|  		|
* 			    	+ve i/p	|
*							-ve i/p
* VCVS gain:
Egain 4 0 2 3 1000
Ebuffer 1 0 5 0 1
* Redundant connection:
Iopen1 2 0 0A
Iopen2 3 0 0A
* Circuit componants:
R1 4 5 1K
C1 5 0 159.15n
.ENDS opamp
.PROBE
.OP
.END
